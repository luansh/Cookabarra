/*-------------------------------------------------------------------------
// Module:  mem
// File:    mem.v
// Author:  shawn Liu
// E-mail:  shawn110285@gmail.com
// Description: LSU
//              (1) handle the load and store instruction
//              (2) process the exception
--------------------------------------------------------------------------*/

`include "defines.v"

module mem(

    input wire n_rst_i,

    /*-- signals from exu-----*/
    input wire[`RegBus] exception_i,       // exception type
    input wire[`RegBus] pc_i,       // the pc when exception happened
    input wire[`RegBus] ins_i,            // the instruction caused the exception

    input wire rd_we_i,
    input wire[`RegAddrBus] rd_wa_i,
    input wire[`RegBus] rd_wd_i,

    input wire[`AluOpBus] uop_i,         //uop_code, to determine it is a load or a store
    input wire[`RegBus] mem_addr_i,
    input wire[`RegBus] mem_wdata_i,

    /*-- signals to access the external memory -----*/
    output reg[`RegBus] mem_a_o,
    output wire mem_we_o,
    output reg[3:0] mem_sel_o,          //the selector for bytes operation
    output reg[`RegBus] mem_data_o,
    output reg mem_ce_o,
    input wire[`RegBus] mem_data_i,        //the read result from memroy

    input wire csr_we_i,
    input wire[`RegBus] csr_waddr_i,
    input wire[`RegBus] csr_wdata_i,

    /*-- signals from write back for data dependance detection -----*/
    input wire wb_csr_we_i,
    input wire[`RegBus] wb_csr_waddr_i,
    input wire[`RegBus] wb_csr_wdata_i,

    /*-- pass down to mem_wb stage -----*/
    output reg rd_we_o,
    output reg[`RegAddrBus] rd_a_o,
    output reg[`RegBus] rd_wd_o,

    output reg csr_we_o,
    output reg[`RegBus] csr_waddr_o,
    output reg[`RegBus] csr_wdata_o,

    /*------- signals to control ----------*/
    output wire stall_req_o,
    output reg[`RegBus] exception_o,
    output reg[`RegBus] pc_o,
    output reg[`RegBus] ins_o

);

    reg mem_we;
    reg mem_re;

    reg addr_align_halfword;
    reg addr_align_word;

    reg load_operation;
    reg store_operation;

    reg load_addr_align_exception;
    reg store_addr_align_exception;

    assign load_operation = ( (uop_i == `UOP_CODE_LH) || (uop_i == `UOP_CODE_LHU) ||(uop_i == `UOP_CODE_LW) ) ? 1'b1 : 1'b0;

    assign store_operation = ( (uop_i == `UOP_CODE_SH) ||(uop_i == `UOP_CODE_SW) ) ? 1'b1 : 1'b0;


    assign addr_align_halfword =(   ( (uop_i == `UOP_CODE_SH) || (uop_i == `UOP_CODE_LH) || (uop_i == `UOP_CODE_LHU) )
                                 && (mem_addr_i[0] == 1'b0) ) ? 1'b1 : 1'b0;

    assign addr_align_word =(   ( (uop_i == `UOP_CODE_SW) || (uop_i == `UOP_CODE_LW) )
                             && (mem_addr_i[1:0] == 2'b00 ) ) ? 1'b1 : 1'b0;

    assign load_addr_align_exception = (~ (addr_align_halfword || addr_align_word)) & load_operation;
    assign store_addr_align_exception = (~ (addr_align_halfword || addr_align_word)) & store_operation;

    // to ctrl module
    //exception ={ misaligned_load, misaligned_store, illegal_inst, misaligned_inst, ebreak, ecall, mret}
    assign exception_o = {25'b0, load_addr_align_exception, store_addr_align_exception, exception_i[4:0]};

    // to the next stage
    assign pc_o = pc_i;
    assign ins_o = ins_i;

    assign csr_we_o = csr_we_i;
    assign csr_waddr_o = csr_waddr_i;
    assign csr_wdata_o = csr_wdata_i;

    assign rd_we_o = rd_we_i;
    assign rd_a_o = rd_wa_i;
    assign rd_wd_o = rd_wd_i;

    assign mem_we = ( (uop_i == `UOP_CODE_SB) || (uop_i == `UOP_CODE_SH)
                    ||(uop_i == `UOP_CODE_SW) ) ? 1'b1 : 1'b0;

    assign mem_re = ( (uop_i == `UOP_CODE_LB) || (uop_i == `UOP_CODE_LBU)
	                ||(uop_i == `UOP_CODE_LH) || (uop_i == `UOP_CODE_LHU)
			   	    ||(uop_i == `UOP_CODE_LW) ) ? 1'b1 : 1'b0;

    assign mem_we_o = mem_we & (~(|exception_o));  // if exeception happened, give up the store operation on the ram
    assign mem_ce_o = mem_we_o | mem_re;
    assign mem_a_o = mem_addr_i;

    assign stall_req_o = 0;

    always @ (*) begin
        if (n_rst_i == `RstEnable) begin
			//operation on RAM
            mem_a_o = `ZeroWord;
            mem_we = `WriteDisable;
            mem_sel_o = 4'b0000;
            mem_data_o = `ZeroWord;
            mem_ce_o = `ChipDisable;

            //GPR
            rd_a_o = `NOPRegAddress;
            rd_we_o = `WriteDisable;
            rd_wd_o = `ZeroWord;

			//CSR
            csr_we_o = `WriteDisable;
            csr_waddr_o = `ZeroWord;
            csr_wdata_o = `ZeroWord;

            exception_o = `ZeroWord;
            pc_o = `ZeroWord;
            ins_o = `NOP_INST;
        end else begin
            mem_sel_o = 4'b1111;
            case (uop_i)
                `UOP_CODE_LB:     begin
                    case (mem_addr_i[1:0])
                        2'b00:  begin
                            rd_wd_o = {{24{mem_data_i[7]}},mem_data_i[7:0]};
                            mem_sel_o = 4'b1000;
                        end
                        2'b01:  begin
                            rd_wd_o = {{24{mem_data_i[15]}},mem_data_i[15:8]};
                            mem_sel_o = 4'b0100;
                        end
                        2'b10:  begin
                            rd_wd_o = {{24{mem_data_i[23]}},mem_data_i[23:16]};
                            mem_sel_o = 4'b0010;
                        end
                        2'b11:  begin
                            rd_wd_o = {{24{mem_data_i[31]}},mem_data_i[31:24]};
                            mem_sel_o = 4'b0001;
                        end
                        default:    begin
                            rd_wd_o = `ZeroWord;
                        end
                    endcase
                end

                `UOP_CODE_LBU:        begin
                    case (mem_addr_i[1:0])
                        2'b00:  begin
                            rd_wd_o = {{24{1'b0}},mem_data_i[7:0]};
                            mem_sel_o = 4'b1000;
                        end
                        2'b01:  begin
                            rd_wd_o = {{24{1'b0}},mem_data_i[15:8]};
                            mem_sel_o = 4'b0100;
                        end
                        2'b10:  begin
                            rd_wd_o = {{24{1'b0}},mem_data_i[23:16]};
                            mem_sel_o = 4'b0010;
                        end
                        2'b11:  begin
                            rd_wd_o = {{24{1'b0}},mem_data_i[31:24]};
                            mem_sel_o = 4'b0001;
                        end
                        default:    begin
                            rd_wd_o = `ZeroWord;
                        end
                    endcase
                end

                `UOP_CODE_LH:     begin
                    case (mem_addr_i[1:0])
                        2'b00:  begin
                            rd_wd_o = {{16{mem_data_i[15]}},mem_data_i[15:0]};
                            mem_sel_o = 4'b1100;
                        end
                        2'b10:  begin
                            rd_wd_o = {{16{mem_data_i[31]}},mem_data_i[31:16]};
                            mem_sel_o = 4'b0011;
                        end
                        default:    begin
                            rd_wd_o = `ZeroWord;
                        end
                    endcase
                end

                `UOP_CODE_LHU:        begin
                    case (mem_addr_i[1:0])
                        2'b00:  begin
                            rd_wd_o = {{16{1'b0}},mem_data_i[15:0]};
                            mem_sel_o = 4'b1100;
                        end
                        2'b10:  begin
                            rd_wd_o = {{16{1'b0}},mem_data_i[31:16]};
                            mem_sel_o = 4'b0011;
                        end
                        default:    begin
                            rd_wd_o = `ZeroWord;
                        end
                    endcase
                end

                `UOP_CODE_LW:     begin
                    rd_wd_o = mem_data_i;
                    mem_sel_o = 4'b1111;
                end

                `UOP_CODE_SB:     begin
                    mem_data_o = {mem_wdata_i[7:0],mem_wdata_i[7:0],mem_wdata_i[7:0],mem_wdata_i[7:0]};
                    case (mem_addr_i[1:0])
                        2'b00:  begin
                            mem_sel_o = 4'b0001;
                        end
                        2'b01:  begin
                            mem_sel_o = 4'b0010;
                        end
                        2'b10:  begin
                            mem_sel_o = 4'b0100;
                        end
                        2'b11:  begin
                            mem_sel_o = 4'b1000;
                        end
                        default:    begin
                            mem_sel_o = 4'b0000;
                        end
                    endcase
                end

                `UOP_CODE_SH:     begin
                    mem_data_o = {mem_wdata_i[15:0],mem_wdata_i[15:0]};
                    case (mem_addr_i[1:0])
                        2'b00:  begin
                            mem_sel_o = 4'b0011;
                        end
                        2'b10:  begin
                            mem_sel_o = 4'b1100;
                        end
                        default:    begin
                            mem_sel_o = 4'b0000;
                        end
                    endcase
                end

                `UOP_CODE_SW:  begin
                    // check the address align with 4 bytes
                    mem_data_o = mem_wdata_i;
                    mem_sel_o = 4'b1111;
                end

                default:  begin
                    //nothing to do
                end
            endcase
        end    //if
    end   //always
endmodule



